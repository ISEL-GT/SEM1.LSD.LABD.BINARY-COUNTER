library ieee;
use ieee.std_logic_1164.all;


-- Entity for counter with control signals
entity binary_counter is

end binary_counter;